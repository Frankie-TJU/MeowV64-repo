../../../build/meowv64.rocket.MeowV64FPGAConfig/meowv64.rocket.MeowV64FPGAConfig.v